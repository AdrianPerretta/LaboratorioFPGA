-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Oct 19 23:50:27 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maquinaestado IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z0 : OUT STD_LOGIC;
        z1 : OUT STD_LOGIC;
        z2 : OUT STD_LOGIC;
        z3 : OUT STD_LOGIC
    );
END maquinaestado;

ARCHITECTURE BEHAVIOR OF maquinaestado IS
    TYPE type_fstate IS (A,C,D,E,B,F,G);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A;
            z0 <= '0';
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
        ELSE
            z0 <= '0';
            z1 <= '0';
            z2 <= '0';
            z3 <= '0';
            CASE fstate IS
                WHEN A =>
                    IF ((x = '0')) THEN
                        reg_fstate <= C;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= D;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A;
                    END IF;

                    z0 <= '0';

                    z1 <= '0';

                    z2 <= '0';

                    z3 <= '0';
                WHEN C =>
                    reg_fstate <= B;

                    z0 <= '0';

                    z1 <= '1';

                    z2 <= '1';

                    z3 <= '0';
                WHEN D =>
                    reg_fstate <= E;

                    z0 <= '0';

                    z1 <= '0';

                    z2 <= '0';

                    z3 <= '1';
                WHEN E =>
                    reg_fstate <= B;

                    z0 <= '0';

                    z1 <= '0';

                    z2 <= '1';

                    z3 <= '1';
                WHEN B =>
                    IF ((x = '1')) THEN
                        reg_fstate <= G;
                    ELSIF ((x = '0')) THEN
                        reg_fstate <= F;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B;
                    END IF;

                    z0 <= '1';

                    z1 <= '1';

                    z2 <= '1';

                    z3 <= '1';
                WHEN F =>
                    reg_fstate <= A;

                    z0 <= '1';

                    z1 <= '0';

                    z2 <= '0';

                    z3 <= '1';
                WHEN G =>
                    reg_fstate <= A;

                    z0 <= '0';

                    z1 <= '1';

                    z2 <= '1';

                    z3 <= '1';
                WHEN OTHERS => 
                    z0 <= 'X';
                    z1 <= 'X';
                    z2 <= 'X';
                    z3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
