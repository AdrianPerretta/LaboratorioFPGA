library verilog;
use verilog.vl_types.all;
entity multModuloCa2_vlg_vec_tst is
end multModuloCa2_vlg_vec_tst;
