-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Oct 31 14:23:34 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mult2bitscs IS 
	PORT
	(
		B0 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		CLEAR :  IN  STD_LOGIC;
		R3 :  OUT  STD_LOGIC;
		R2 :  OUT  STD_LOGIC;
		R1 :  OUT  STD_LOGIC;
		R0 :  OUT  STD_LOGIC;
		BANDERA_CEROS :  OUT  STD_LOGIC;
		BANDERA_SIGNO :  OUT  STD_LOGIC
	);
END mult2bitscs;

ARCHITECTURE bdf_type OF mult2bitscs IS 

COMPONENT fulladder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 COUT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	DFF_inst16 :  STD_LOGIC;
SIGNAL	DFF_inst17 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;


BEGIN 
R3 <= SYNTHESIZED_WIRE_45;
R2 <= DFF_inst16;
R1 <= DFF_inst17;
R0 <= DFF_inst18;
BANDERA_SIGNO <= SYNTHESIZED_WIRE_45;
SYNTHESIZED_WIRE_40 <= '0';
SYNTHESIZED_WIRE_42 <= '1';
SYNTHESIZED_WIRE_43 <= '1';
SYNTHESIZED_WIRE_21 <= '0';
SYNTHESIZED_WIRE_36 <= '1';





SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38;


b2v_inst12 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_40,
		 CIN => SYNTHESIZED_WIRE_2,
		 S => SYNTHESIZED_WIRE_32,
		 COUT => SYNTHESIZED_WIRE_27);


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_41;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_42)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_45 <= '0';
ELSIF (SYNTHESIZED_WIRE_42 = '0') THEN
	SYNTHESIZED_WIRE_45 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_45 <= SYNTHESIZED_WIRE_4;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_42)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst16 <= '0';
ELSIF (SYNTHESIZED_WIRE_42 = '0') THEN
	DFF_inst16 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst16 <= SYNTHESIZED_WIRE_6;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_42)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst17 <= '0';
ELSIF (SYNTHESIZED_WIRE_42 = '0') THEN
	DFF_inst17 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst17 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_42)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_42 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst18 <= SYNTHESIZED_WIRE_10;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_43)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_37 <= '0';
ELSIF (SYNTHESIZED_WIRE_43 = '0') THEN
	SYNTHESIZED_WIRE_37 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_37 <= A1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_10 <= SYNTHESIZED_WIRE_44 AND SYNTHESIZED_WIRE_38;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_43)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_44 <= '0';
ELSIF (SYNTHESIZED_WIRE_43 = '0') THEN
	SYNTHESIZED_WIRE_44 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_44 <= A0;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_43)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_38 <= '0';
ELSIF (SYNTHESIZED_WIRE_43 = '0') THEN
	SYNTHESIZED_WIRE_38 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_38 <= B0;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_43)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_41 <= '0';
ELSIF (SYNTHESIZED_WIRE_43 = '0') THEN
	SYNTHESIZED_WIRE_41 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_41 <= B1;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38;



b2v_inst26 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_16,
		 B => SYNTHESIZED_WIRE_17,
		 CIN => SYNTHESIZED_WIRE_18,
		 S => SYNTHESIZED_WIRE_6,
		 COUT => SYNTHESIZED_WIRE_24);


b2v_inst27 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_19,
		 B => SYNTHESIZED_WIRE_20,
		 CIN => SYNTHESIZED_WIRE_21,
		 S => SYNTHESIZED_WIRE_8,
		 COUT => SYNTHESIZED_WIRE_18);


b2v_inst28 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_22,
		 B => SYNTHESIZED_WIRE_23,
		 CIN => SYNTHESIZED_WIRE_24,
		 S => SYNTHESIZED_WIRE_4);


b2v_inst29 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_40,
		 CIN => SYNTHESIZED_WIRE_27,
		 S => SYNTHESIZED_WIRE_3);


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38;


BANDERA_CEROS <= SYNTHESIZED_WIRE_28 AND SYNTHESIZED_WIRE_29 AND SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_28 <= NOT(SYNTHESIZED_WIRE_45);



SYNTHESIZED_WIRE_29 <= NOT(DFF_inst16);



SYNTHESIZED_WIRE_30 <= NOT(DFF_inst17);



SYNTHESIZED_WIRE_31 <= NOT(DFF_inst18);



SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_32 AND SYNTHESIZED_WIRE_41;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_41;



b2v_inst7 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_34,
		 B => SYNTHESIZED_WIRE_40,
		 CIN => SYNTHESIZED_WIRE_36,
		 S => SYNTHESIZED_WIRE_33,
		 COUT => SYNTHESIZED_WIRE_2);


SYNTHESIZED_WIRE_34 <= NOT(SYNTHESIZED_WIRE_44);



SYNTHESIZED_WIRE_39 <= NOT(SYNTHESIZED_WIRE_37);



END bdf_type;