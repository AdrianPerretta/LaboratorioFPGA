library verilog;
use verilog.vl_types.all;
entity maquinaestado_vlg_check_tst is
    port(
        z0              : in     vl_logic;
        z1              : in     vl_logic;
        z2              : in     vl_logic;
        z3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end maquinaestado_vlg_check_tst;
