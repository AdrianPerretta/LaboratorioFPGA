library verilog;
use verilog.vl_types.all;
entity maquinaestado_vlg_vec_tst is
end maquinaestado_vlg_vec_tst;
