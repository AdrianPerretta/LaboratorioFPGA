-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Wed Oct 29 20:54:56 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY i2c IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        Hab_dir : OUT STD_LOGIC;
        Hab_dato : OUT STD_LOGIC;
        acknowledge : OUT STD_LOGIC
    );
END i2c;

ARCHITECTURE BEHAVIOR OF i2c IS
    TYPE type_fstate IS (Oscioso,Guardar_dir,ROW,ACK_Estado,Guardar_Dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,fin_dir,fin_dato,soy)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Oscioso;
            Hab_dir <= '0';
            Hab_dato <= '0';
            acknowledge <= '0';
        ELSE
            Hab_dir <= '0';
            Hab_dato <= '0';
            acknowledge <= '0';
            CASE fstate IS
                WHEN Oscioso =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= Oscioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Oscioso;
                    END IF;

                    acknowledge <= '0';

                    Hab_dir <= '0';

                    Hab_dato <= '0';
                WHEN Guardar_dir =>
                    IF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= ROW;
                    ELSIF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guardar_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_dir;
                    END IF;

                    acknowledge <= '0';

                    Hab_dir <= '1';

                    Hab_dato <= '0';
                WHEN ROW =>
                    reg_fstate <= ACK_Estado;

                    acknowledge <= '0';

                    Hab_dir <= '0';

                    Hab_dato <= '0';
                WHEN ACK_Estado =>
                    reg_fstate <= Guardar_Dato;

                    acknowledge <= '1';

                    Hab_dir <= '0';

                    Hab_dato <= '0';
                WHEN Guardar_Dato =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= Oscioso;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= Guardar_Dato;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guardar_Dato;
                    END IF;

                    acknowledge <= '0';

                    Hab_dir <= '0';

                    Hab_dato <= '1';
                WHEN OTHERS => 
                    Hab_dir <= 'X';
                    Hab_dato <= 'X';
                    acknowledge <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
