library verilog;
use verilog.vl_types.all;
entity mult2bits_vlg_vec_tst is
end mult2bits_vlg_vec_tst;
