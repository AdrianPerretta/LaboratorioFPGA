-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Tue Oct 28 23:05:24 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mult2bitscs IS 
	PORT
	(
		B0 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		CLEAR :  IN  STD_LOGIC;
		R3 :  OUT  STD_LOGIC;
		R2 :  OUT  STD_LOGIC;
		R1 :  OUT  STD_LOGIC;
		R0 :  OUT  STD_LOGIC;
		BANDERA_CEROS :  OUT  STD_LOGIC;
		BANDERA_SIGNO :  OUT  STD_LOGIC
	);
END mult2bitscs;

ARCHITECTURE bdf_type OF mult2bitscs IS 

COMPONENT fulladder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 COUT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	DFF_inst16 :  STD_LOGIC;
SIGNAL	DFF_inst17 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;


BEGIN 
R3 <= SYNTHESIZED_WIRE_41;
R2 <= DFF_inst16;
R1 <= DFF_inst17;
R0 <= DFF_inst18;
BANDERA_SIGNO <= SYNTHESIZED_WIRE_41;
SYNTHESIZED_WIRE_36 <= '0';
SYNTHESIZED_WIRE_37 <= '1';
SYNTHESIZED_WIRE_38 <= '1';
SYNTHESIZED_WIRE_22 <= '0';
SYNTHESIZED_WIRE_33 <= '1';



SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1;




SYNTHESIZED_WIRE_18 <= SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35;


b2v_inst12 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_2,
		 B => SYNTHESIZED_WIRE_36,
		 CIN => SYNTHESIZED_WIRE_4,
		 S => SYNTHESIZED_WIRE_29);


SYNTHESIZED_WIRE_23 <= NOT(SYNTHESIZED_WIRE_34);



PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_37)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_41 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	SYNTHESIZED_WIRE_41 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_41 <= SYNTHESIZED_WIRE_5;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_37)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst16 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst16 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst16 <= SYNTHESIZED_WIRE_7;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_37)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst17 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst17 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst17 <= SYNTHESIZED_WIRE_9;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_37)
BEGIN
IF (CLEAR = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_37 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst18 <= SYNTHESIZED_WIRE_11;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_38)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_34 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	SYNTHESIZED_WIRE_34 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_34 <= A1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_11 <= SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_35;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_38)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_39 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	SYNTHESIZED_WIRE_39 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_39 <= A0;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_38)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_35 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	SYNTHESIZED_WIRE_35 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_35 <= B0;
END IF;
END PROCESS;


PROCESS(CLK,CLEAR,SYNTHESIZED_WIRE_38)
BEGIN
IF (CLEAR = '0') THEN
	SYNTHESIZED_WIRE_40 <= '0';
ELSIF (SYNTHESIZED_WIRE_38 = '0') THEN
	SYNTHESIZED_WIRE_40 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_40 <= B1;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_24 <= NOT(SYNTHESIZED_WIRE_40);




b2v_inst26 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_17,
		 B => SYNTHESIZED_WIRE_18,
		 CIN => SYNTHESIZED_WIRE_19,
		 S => SYNTHESIZED_WIRE_7);


b2v_inst27 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_20,
		 B => SYNTHESIZED_WIRE_21,
		 CIN => SYNTHESIZED_WIRE_22,
		 S => SYNTHESIZED_WIRE_9,
		 COUT => SYNTHESIZED_WIRE_19);


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_23 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35 AND SYNTHESIZED_WIRE_24;


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35;


BANDERA_CEROS <= SYNTHESIZED_WIRE_25 AND SYNTHESIZED_WIRE_26 AND SYNTHESIZED_WIRE_27 AND SYNTHESIZED_WIRE_28;


SYNTHESIZED_WIRE_25 <= NOT(SYNTHESIZED_WIRE_41);



SYNTHESIZED_WIRE_26 <= NOT(DFF_inst16);



SYNTHESIZED_WIRE_27 <= NOT(DFF_inst17);



SYNTHESIZED_WIRE_28 <= NOT(DFF_inst18);



SYNTHESIZED_WIRE_17 <= SYNTHESIZED_WIRE_29 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_20 <= SYNTHESIZED_WIRE_30 AND SYNTHESIZED_WIRE_40;



b2v_inst7 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_31,
		 B => SYNTHESIZED_WIRE_36,
		 CIN => SYNTHESIZED_WIRE_33,
		 S => SYNTHESIZED_WIRE_30,
		 COUT => SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_31 <= NOT(SYNTHESIZED_WIRE_39);



SYNTHESIZED_WIRE_2 <= NOT(SYNTHESIZED_WIRE_34);



END bdf_type;