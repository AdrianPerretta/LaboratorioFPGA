-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Fri Oct 24 12:02:00 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY mult2bitscs IS 
	PORT
	(
		B0 :  IN  STD_LOGIC;
		A0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		R3 :  OUT  STD_LOGIC;
		R2 :  OUT  STD_LOGIC;
		R1 :  OUT  STD_LOGIC;
		R0 :  OUT  STD_LOGIC;
		BANDERA_CEROS :  OUT  STD_LOGIC;
		BANDERA_SIGNO :  OUT  STD_LOGIC
	);
END mult2bitscs;

ARCHITECTURE bdf_type OF mult2bitscs IS 

COMPONENT fulladder
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 CIN : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 COUT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_45 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_46 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_47 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_34 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_35 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_36 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_49 :  STD_LOGIC;
SIGNAL	DFF_inst16 :  STD_LOGIC;
SIGNAL	DFF_inst17 :  STD_LOGIC;
SIGNAL	DFF_inst18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;


BEGIN 
R3 <= SYNTHESIZED_WIRE_49;
R2 <= DFF_inst16;
R1 <= DFF_inst17;
R0 <= DFF_inst18;
BANDERA_SIGNO <= SYNTHESIZED_WIRE_49;
SYNTHESIZED_WIRE_44 <= '0';
SYNTHESIZED_WIRE_45 <= '1';
SYNTHESIZED_WIRE_46 <= '1';
SYNTHESIZED_WIRE_30 <= '0';
SYNTHESIZED_WIRE_41 <= '1';



SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_0 OR SYNTHESIZED_WIRE_1;




SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


b2v_inst12 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_2,
		 B => SYNTHESIZED_WIRE_44,
		 CIN => SYNTHESIZED_WIRE_4,
		 S => SYNTHESIZED_WIRE_37);


SYNTHESIZED_WIRE_31 <= NOT(SYNTHESIZED_WIRE_42);



PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_49 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	SYNTHESIZED_WIRE_49 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_49 <= SYNTHESIZED_WIRE_6;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst16 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst16 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst16 <= SYNTHESIZED_WIRE_9;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst17 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst17 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst17 <= SYNTHESIZED_WIRE_12;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_45,SYNTHESIZED_WIRE_45)
BEGIN
IF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst18 <= '0';
ELSIF (SYNTHESIZED_WIRE_45 = '0') THEN
	DFF_inst18 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	DFF_inst18 <= SYNTHESIZED_WIRE_15;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_46,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_42 <= '0';
ELSIF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_42 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_42 <= A1;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_15 <= SYNTHESIZED_WIRE_47 AND SYNTHESIZED_WIRE_43;


PROCESS(CLK,SYNTHESIZED_WIRE_46,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '0';
ELSIF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_47 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_47 <= A0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_46,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '0';
ELSIF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_43 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_43 <= B0;
END IF;
END PROCESS;


PROCESS(CLK,SYNTHESIZED_WIRE_46,SYNTHESIZED_WIRE_46)
BEGIN
IF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_48 <= '0';
ELSIF (SYNTHESIZED_WIRE_46 = '0') THEN
	SYNTHESIZED_WIRE_48 <= '1';
ELSIF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_48 <= B1;
END IF;
END PROCESS;



SYNTHESIZED_WIRE_32 <= NOT(SYNTHESIZED_WIRE_48);




b2v_inst26 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_25,
		 B => SYNTHESIZED_WIRE_26,
		 CIN => SYNTHESIZED_WIRE_27,
		 S => SYNTHESIZED_WIRE_9);


b2v_inst27 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_28,
		 B => SYNTHESIZED_WIRE_29,
		 CIN => SYNTHESIZED_WIRE_30,
		 S => SYNTHESIZED_WIRE_12,
		 COUT => SYNTHESIZED_WIRE_27);


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_47 AND SYNTHESIZED_WIRE_31 AND SYNTHESIZED_WIRE_48;


SYNTHESIZED_WIRE_0 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_29 <= SYNTHESIZED_WIRE_42 AND SYNTHESIZED_WIRE_43;


BANDERA_CEROS <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_34 AND SYNTHESIZED_WIRE_35 AND SYNTHESIZED_WIRE_36;


SYNTHESIZED_WIRE_33 <= NOT(SYNTHESIZED_WIRE_49);



SYNTHESIZED_WIRE_34 <= NOT(DFF_inst16);



SYNTHESIZED_WIRE_35 <= NOT(DFF_inst17);



SYNTHESIZED_WIRE_36 <= NOT(DFF_inst18);



SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_48;


SYNTHESIZED_WIRE_28 <= SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_48;



b2v_inst7 : fulladder
PORT MAP(A => SYNTHESIZED_WIRE_39,
		 B => SYNTHESIZED_WIRE_44,
		 CIN => SYNTHESIZED_WIRE_41,
		 S => SYNTHESIZED_WIRE_38,
		 COUT => SYNTHESIZED_WIRE_4);


SYNTHESIZED_WIRE_39 <= NOT(SYNTHESIZED_WIRE_47);



SYNTHESIZED_WIRE_2 <= NOT(SYNTHESIZED_WIRE_42);



END bdf_type;