library verilog;
use verilog.vl_types.all;
entity i2cEsquematico_vlg_vec_tst is
end i2cEsquematico_vlg_vec_tst;
