library verilog;
use verilog.vl_types.all;
entity mult2bitscs_vlg_vec_tst is
end mult2bitscs_vlg_vec_tst;
